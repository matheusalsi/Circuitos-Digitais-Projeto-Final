library verilog;
use verilog.vl_types.all;
entity mod3_bcd_vlg_vec_tst is
end mod3_bcd_vlg_vec_tst;
