library verilog;
use verilog.vl_types.all;
entity sixbit_inc_register_vlg_vec_tst is
end sixbit_inc_register_vlg_vec_tst;
