library verilog;
use verilog.vl_types.all;
entity sixbit_to_bcd_vlg_vec_tst is
end sixbit_to_bcd_vlg_vec_tst;
