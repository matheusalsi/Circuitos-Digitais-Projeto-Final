library verilog;
use verilog.vl_types.all;
entity cronometer_control_vlg_vec_tst is
end cronometer_control_vlg_vec_tst;
