library verilog;
use verilog.vl_types.all;
entity trabalho_final_vlg_vec_tst is
end trabalho_final_vlg_vec_tst;
