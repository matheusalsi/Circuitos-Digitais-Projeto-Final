library verilog;
use verilog.vl_types.all;
entity cr_counter_vlg_vec_tst is
end cr_counter_vlg_vec_tst;
