library verilog;
use verilog.vl_types.all;
entity mod60_counter_vlg_vec_tst is
end mod60_counter_vlg_vec_tst;
